module moduleNamePlaceholder (
);
    
endmodule